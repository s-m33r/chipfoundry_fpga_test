VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 309.440 500.000 310.040 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 496.000 261.190 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 336.640 500.000 337.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 479.440 500.000 480.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 496.000 132.390 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 34.040 500.000 34.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 496.000 71.210 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 496.000 174.250 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 496.000 335.250 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 326.440 500.000 327.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 37.440 500.000 38.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 496.000 180.690 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 496.000 103.410 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 496.000 148.490 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 496.000 380.330 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.840 500.000 313.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 391.040 500.000 391.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 496.000 460.830 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END prog_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 494.280 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 494.280 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 494.280 334.690 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 487.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 494.280 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 494.280 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 494.280 337.990 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.760 494.230 487.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.530 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 0.550 495.720 67.430 496.810 ;
        RECT 68.270 495.720 70.650 496.810 ;
        RECT 71.490 495.720 102.850 496.810 ;
        RECT 103.690 495.720 131.830 496.810 ;
        RECT 132.670 495.720 147.930 496.810 ;
        RECT 148.770 495.720 173.690 496.810 ;
        RECT 174.530 495.720 180.130 496.810 ;
        RECT 180.970 495.720 260.630 496.810 ;
        RECT 261.470 495.720 334.690 496.810 ;
        RECT 335.530 495.720 350.790 496.810 ;
        RECT 351.630 495.720 376.550 496.810 ;
        RECT 377.390 495.720 379.770 496.810 ;
        RECT 380.610 495.720 460.270 496.810 ;
        RECT 461.110 495.720 492.570 496.810 ;
        RECT 0.550 4.280 492.570 495.720 ;
        RECT 0.650 4.000 3.030 4.280 ;
        RECT 3.870 4.000 6.250 4.280 ;
        RECT 7.090 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 231.650 4.280 ;
        RECT 232.490 4.000 263.850 4.280 ;
        RECT 264.690 4.000 308.930 4.280 ;
        RECT 309.770 4.000 315.370 4.280 ;
        RECT 316.210 4.000 321.810 4.280 ;
        RECT 322.650 4.000 360.450 4.280 ;
        RECT 361.290 4.000 466.710 4.280 ;
        RECT 467.550 4.000 476.370 4.280 ;
        RECT 477.210 4.000 492.570 4.280 ;
      LAYER met3 ;
        RECT 0.525 483.840 496.000 487.045 ;
        RECT 0.525 482.440 495.600 483.840 ;
        RECT 0.525 480.440 496.000 482.440 ;
        RECT 0.525 479.040 495.600 480.440 ;
        RECT 0.525 466.840 496.000 479.040 ;
        RECT 4.400 465.440 496.000 466.840 ;
        RECT 0.525 463.440 496.000 465.440 ;
        RECT 4.400 462.040 496.000 463.440 ;
        RECT 0.525 405.640 496.000 462.040 ;
        RECT 0.525 404.240 495.600 405.640 ;
        RECT 0.525 392.040 496.000 404.240 ;
        RECT 0.525 390.640 495.600 392.040 ;
        RECT 0.525 385.240 496.000 390.640 ;
        RECT 4.400 383.840 496.000 385.240 ;
        RECT 0.525 344.440 496.000 383.840 ;
        RECT 0.525 343.040 495.600 344.440 ;
        RECT 0.525 341.040 496.000 343.040 ;
        RECT 0.525 339.640 495.600 341.040 ;
        RECT 0.525 337.640 496.000 339.640 ;
        RECT 0.525 336.240 495.600 337.640 ;
        RECT 0.525 327.440 496.000 336.240 ;
        RECT 0.525 326.040 495.600 327.440 ;
        RECT 0.525 313.840 496.000 326.040 ;
        RECT 0.525 312.440 495.600 313.840 ;
        RECT 0.525 310.440 496.000 312.440 ;
        RECT 0.525 309.040 495.600 310.440 ;
        RECT 0.525 266.240 496.000 309.040 ;
        RECT 0.525 264.840 495.600 266.240 ;
        RECT 0.525 218.640 496.000 264.840 ;
        RECT 0.525 217.240 495.600 218.640 ;
        RECT 0.525 208.440 496.000 217.240 ;
        RECT 4.400 207.040 496.000 208.440 ;
        RECT 0.525 184.640 496.000 207.040 ;
        RECT 4.400 183.240 496.000 184.640 ;
        RECT 0.525 147.240 496.000 183.240 ;
        RECT 4.400 145.840 496.000 147.240 ;
        RECT 0.525 123.440 496.000 145.840 ;
        RECT 4.400 122.040 496.000 123.440 ;
        RECT 0.525 103.040 496.000 122.040 ;
        RECT 0.525 101.640 495.600 103.040 ;
        RECT 0.525 96.240 496.000 101.640 ;
        RECT 0.525 94.840 495.600 96.240 ;
        RECT 0.525 52.040 496.000 94.840 ;
        RECT 0.525 50.640 495.600 52.040 ;
        RECT 0.525 45.240 496.000 50.640 ;
        RECT 0.525 43.840 495.600 45.240 ;
        RECT 0.525 41.840 496.000 43.840 ;
        RECT 0.525 40.440 495.600 41.840 ;
        RECT 0.525 38.440 496.000 40.440 ;
        RECT 0.525 37.040 495.600 38.440 ;
        RECT 0.525 35.040 496.000 37.040 ;
        RECT 0.525 33.640 495.600 35.040 ;
        RECT 0.525 10.715 496.000 33.640 ;
  END
END fpga_top
END LIBRARY

