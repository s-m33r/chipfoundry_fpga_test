//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Nov 26 15:27:55 2025
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(clk,
                IO_ISOL_N,
                prog_clk,
                Test_en,
                gfpga_pad_EMBEDDED_IO_HD_SOC_IN,
                gfpga_pad_EMBEDDED_IO_HD_SOC_OUT,
                gfpga_pad_EMBEDDED_IO_HD_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GPIN PORTS -----
input [0:23] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
//----- GPOUT PORTS -----
output [0:23] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
//----- GPOUT PORTS -----
output [0:23] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:19] cbx_1__0__0_chanx_left_out;
wire [0:19] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:19] cbx_1__0__1_chanx_left_out;
wire [0:19] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:19] cbx_1__1__0_chanx_left_out;
wire [0:19] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:19] cbx_1__1__1_chanx_left_out;
wire [0:19] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:19] cbx_1__2__0_chanx_left_out;
wire [0:19] cbx_1__2__0_chanx_right_out;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:19] cbx_1__2__1_chanx_left_out;
wire [0:19] cbx_1__2__1_chanx_right_out;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:19] cby_0__1__0_chany_bottom_out;
wire [0:19] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:19] cby_0__1__1_chany_bottom_out;
wire [0:19] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:19] cby_1__1__0_chany_bottom_out;
wire [0:19] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:19] cby_1__1__1_chany_bottom_out;
wire [0:19] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_2__1__0_ccff_tail;
wire [0:19] cby_2__1__0_chany_bottom_out;
wire [0:19] cby_2__1__0_chany_top_out;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_2__1__1_ccff_tail;
wire [0:19] cby_2__1__1_chany_bottom_out;
wire [0:19] cby_2__1__1_chany_top_out;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_;
wire [0:0] cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_;
wire [0:0] cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_1_out;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_;
wire [0:0] grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_upper;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_lower;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_upper;
wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_0_ccff_tail;
wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_left_left_1_ccff_tail;
wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_0_ccff_tail;
wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_right_right_1_ccff_tail;
wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_0_ccff_tail;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper;
wire [0:0] grid_io_top_top_1_ccff_tail;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:19] sb_0__0__0_chanx_right_out;
wire [0:19] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:19] sb_0__1__0_chanx_right_out;
wire [0:19] sb_0__1__0_chany_bottom_out;
wire [0:19] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:19] sb_0__2__0_chanx_right_out;
wire [0:19] sb_0__2__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:19] sb_1__0__0_chanx_left_out;
wire [0:19] sb_1__0__0_chanx_right_out;
wire [0:19] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:19] sb_1__1__0_chanx_left_out;
wire [0:19] sb_1__1__0_chanx_right_out;
wire [0:19] sb_1__1__0_chany_bottom_out;
wire [0:19] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:19] sb_1__2__0_chanx_left_out;
wire [0:19] sb_1__2__0_chanx_right_out;
wire [0:19] sb_1__2__0_chany_bottom_out;
wire [0:0] sb_2__0__0_ccff_tail;
wire [0:19] sb_2__0__0_chanx_left_out;
wire [0:19] sb_2__0__0_chany_top_out;
wire [0:0] sb_2__1__0_ccff_tail;
wire [0:19] sb_2__1__0_chanx_left_out;
wire [0:19] sb_2__1__0_chany_bottom_out;
wire [0:19] sb_2__1__0_chany_top_out;
wire [0:0] sb_2__2__0_ccff_tail;
wire [0:19] sb_2__2__0_chanx_left_out;
wire [0:19] sb_2__2__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top_top grid_io_top_top_1__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_top_top_1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_0_ccff_tail));

	grid_io_top_top grid_io_top_top_2__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_top_top_1_ccff_tail));

	grid_io_right_right grid_io_right_right_3__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_0_ccff_tail));

	grid_io_right_right grid_io_right_right_3__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.left_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_right_right_1_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_2__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4:12]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4:12]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4:12]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_0_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_1__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13:21]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13:21]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13:21]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_1__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_1__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_2__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_2__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_3__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_3__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_4__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_4__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_5__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_5__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_6__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_6__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_7__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_7__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.top_width_0_height_0_subtile_8__pin_inpad_0_upper(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.top_width_0_height_0_subtile_8__pin_inpad_0_lower(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_tail(grid_io_bottom_bottom_1_ccff_tail));

	grid_io_left_left grid_io_left_left_0__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_0_ccff_tail));

	grid_io_left_left grid_io_left_left_0__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_upper(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_width_0_height_0_subtile_0__pin_inpad_0_lower(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.ccff_tail(grid_io_left_left_1_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.top_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.top_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.right_width_0_height_0_subtile_0__pin_O_12_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.right_width_0_height_0_subtile_0__pin_O_12_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.right_width_0_height_0_subtile_0__pin_O_13_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.right_width_0_height_0_subtile_0__pin_O_13_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.right_width_0_height_0_subtile_0__pin_O_14_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.right_width_0_height_0_subtile_0__pin_O_14_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.right_width_0_height_0_subtile_0__pin_O_15_upper(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.right_width_0_height_0_subtile_0__pin_O_15_lower(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.top_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.top_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.right_width_0_height_0_subtile_0__pin_O_12_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.right_width_0_height_0_subtile_0__pin_O_12_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.right_width_0_height_0_subtile_0__pin_O_13_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.right_width_0_height_0_subtile_0__pin_O_13_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.right_width_0_height_0_subtile_0__pin_O_14_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.right_width_0_height_0_subtile_0__pin_O_14_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.right_width_0_height_0_subtile_0__pin_O_15_upper(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.right_width_0_height_0_subtile_0__pin_O_15_lower(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_0_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_1_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_2__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.top_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.top_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.right_width_0_height_0_subtile_0__pin_O_12_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.right_width_0_height_0_subtile_0__pin_O_12_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.right_width_0_height_0_subtile_0__pin_O_13_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.right_width_0_height_0_subtile_0__pin_O_13_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.right_width_0_height_0_subtile_0__pin_O_14_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.right_width_0_height_0_subtile_0__pin_O_14_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.right_width_0_height_0_subtile_0__pin_O_15_upper(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.right_width_0_height_0_subtile_0__pin_O_15_lower(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_2__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.top_width_0_height_0_subtile_0__pin_O_0_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.top_width_0_height_0_subtile_0__pin_O_1_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.top_width_0_height_0_subtile_0__pin_O_1_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.top_width_0_height_0_subtile_0__pin_O_2_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.top_width_0_height_0_subtile_0__pin_O_2_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.top_width_0_height_0_subtile_0__pin_O_3_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.top_width_0_height_0_subtile_0__pin_O_3_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.top_width_0_height_0_subtile_0__pin_O_4_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.top_width_0_height_0_subtile_0__pin_O_4_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.top_width_0_height_0_subtile_0__pin_O_5_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.top_width_0_height_0_subtile_0__pin_O_5_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.top_width_0_height_0_subtile_0__pin_O_6_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.top_width_0_height_0_subtile_0__pin_O_6_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.top_width_0_height_0_subtile_0__pin_O_7_upper(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.top_width_0_height_0_subtile_0__pin_O_7_lower(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.right_width_0_height_0_subtile_0__pin_O_8_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.right_width_0_height_0_subtile_0__pin_O_8_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.right_width_0_height_0_subtile_0__pin_O_9_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.right_width_0_height_0_subtile_0__pin_O_9_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.right_width_0_height_0_subtile_0__pin_O_10_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.right_width_0_height_0_subtile_0__pin_O_10_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.right_width_0_height_0_subtile_0__pin_O_11_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.right_width_0_height_0_subtile_0__pin_O_11_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.right_width_0_height_0_subtile_0__pin_O_12_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.right_width_0_height_0_subtile_0__pin_O_12_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.right_width_0_height_0_subtile_0__pin_O_13_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.right_width_0_height_0_subtile_0__pin_O_13_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.right_width_0_height_0_subtile_0__pin_O_14_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.right_width_0_height_0_subtile_0__pin_O_14_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.right_width_0_height_0_subtile_0__pin_O_15_upper(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.right_width_0_height_0_subtile_0__pin_O_15_lower(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(grid_clb_3_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.ccff_head(ccff_head),
		.chany_top_out(sb_0__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_left_left_1_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__2_ sb_0__2_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__2__0_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_head(grid_io_top_top_0_ccff_tail),
		.chanx_right_out(sb_0__2__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__2__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__2__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.ccff_head(grid_io_left_left_0_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__2__1_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_upper),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_upper),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.chanx_left_in(cbx_1__2__0_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.ccff_head(grid_clb_3_ccff_tail),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_2__0_ sb_2__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_8__pin_inpad_0_lower),
		.ccff_head(grid_io_bottom_bottom_1_ccff_tail),
		.chany_top_out(sb_2__0__0_chany_top_out[0:19]),
		.chanx_left_out(sb_2__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_2__0__0_ccff_tail));

	sb_2__1_ sb_2__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_lower),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_lower),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.chany_bottom_in(cby_2__1__0_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_2__1__0_chany_top_out[0:19]),
		.chany_bottom_out(sb_2__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_2__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_2__1__0_ccff_tail));

	sb_2__2_ sb_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_2__1__1_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_upper),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_upper),
		.chanx_left_in(cbx_1__2__1_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_lower),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_lower),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_bottom_out(sb_2__2__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_2__2__0_chanx_left_out[0:19]),
		.ccff_tail(sb_2__2__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_2__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_2__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_2__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_2__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__2_ cbx_1__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__2__0_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__2__0_ccff_tail));

	cbx_1__2_ cbx_2__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_2__2__0_chanx_left_out[0:19]),
		.ccff_head(sb_2__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__2__1_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.ccff_tail(cbx_1__2__1_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:19]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__2__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__2__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:19]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:19]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__2__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:19]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_2__1_ cby_2__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_2__1__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_2__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_2__1__0_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_2__1__0_ccff_tail));

	cby_2__1_ cby_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_2__2__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__2__1_ccff_tail),
		.chany_bottom_out(cby_2__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_2__1__1_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_2_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_2__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.ccff_tail(cby_2__1__1_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_1_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




