VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.840 500.000 347.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 496.000 74.430 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 496.000 116.290 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 496.000 77.650 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 241.440 500.000 242.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 496.000 167.810 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 496.000 338.470 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 47.640 500.000 48.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 496.000 190.350 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 496.000 106.630 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 496.000 151.710 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 496.000 357.790 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 136.040 500.000 136.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 54.440 500.000 55.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 496.000 367.450 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 496.000 451.170 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 496.000 454.390 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 496.000 51.890 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 435.240 500.000 435.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 496.000 447.950 500.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 64.640 500.000 65.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END prog_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 43.470 40.560 46.570 459.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.470 40.560 226.570 459.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 403.470 40.560 406.570 459.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 44.250 460.240 47.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 224.250 460.240 227.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 404.250 460.240 407.350 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 62.070 40.560 65.170 459.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 242.070 40.560 245.170 459.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 422.070 40.560 425.170 459.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 62.850 460.240 65.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 242.850 460.240 245.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 39.780 422.850 460.240 425.950 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 39.830 40.715 460.190 459.765 ;
      LAYER li1 ;
        RECT 40.020 40.715 460.000 459.765 ;
      LAYER met1 ;
        RECT 0.530 40.560 491.210 483.100 ;
      LAYER met2 ;
        RECT 0.550 495.720 51.330 496.810 ;
        RECT 52.170 495.720 54.550 496.810 ;
        RECT 55.390 495.720 73.870 496.810 ;
        RECT 74.710 495.720 77.090 496.810 ;
        RECT 77.930 495.720 106.070 496.810 ;
        RECT 106.910 495.720 115.730 496.810 ;
        RECT 116.570 495.720 151.150 496.810 ;
        RECT 151.990 495.720 167.250 496.810 ;
        RECT 168.090 495.720 189.790 496.810 ;
        RECT 190.630 495.720 331.470 496.810 ;
        RECT 332.310 495.720 337.910 496.810 ;
        RECT 338.750 495.720 357.230 496.810 ;
        RECT 358.070 495.720 366.890 496.810 ;
        RECT 367.730 495.720 376.550 496.810 ;
        RECT 377.390 495.720 444.170 496.810 ;
        RECT 445.010 495.720 447.390 496.810 ;
        RECT 448.230 495.720 450.610 496.810 ;
        RECT 451.450 495.720 453.830 496.810 ;
        RECT 454.670 495.720 491.190 496.810 ;
        RECT 0.550 4.280 491.190 495.720 ;
        RECT 0.650 4.000 3.030 4.280 ;
        RECT 3.870 4.000 6.250 4.280 ;
        RECT 7.090 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 151.150 4.280 ;
        RECT 151.990 4.000 283.170 4.280 ;
        RECT 284.010 4.000 292.830 4.280 ;
        RECT 293.670 4.000 315.370 4.280 ;
        RECT 316.210 4.000 331.470 4.280 ;
        RECT 332.310 4.000 347.570 4.280 ;
        RECT 348.410 4.000 447.390 4.280 ;
        RECT 448.230 4.000 491.190 4.280 ;
      LAYER met3 ;
        RECT 0.525 436.240 496.000 459.845 ;
        RECT 0.525 434.840 495.600 436.240 ;
        RECT 0.525 426.040 496.000 434.840 ;
        RECT 4.400 424.640 496.000 426.040 ;
        RECT 0.525 388.640 496.000 424.640 ;
        RECT 0.525 387.240 495.600 388.640 ;
        RECT 0.525 347.840 496.000 387.240 ;
        RECT 0.525 346.440 495.600 347.840 ;
        RECT 0.525 344.440 496.000 346.440 ;
        RECT 0.525 343.040 495.600 344.440 ;
        RECT 0.525 341.040 496.000 343.040 ;
        RECT 0.525 339.640 495.600 341.040 ;
        RECT 0.525 262.840 496.000 339.640 ;
        RECT 4.400 261.440 495.600 262.840 ;
        RECT 0.525 242.440 496.000 261.440 ;
        RECT 4.400 241.040 495.600 242.440 ;
        RECT 0.525 188.040 496.000 241.040 ;
        RECT 0.525 186.640 495.600 188.040 ;
        RECT 0.525 167.640 496.000 186.640 ;
        RECT 4.400 166.240 496.000 167.640 ;
        RECT 0.525 147.240 496.000 166.240 ;
        RECT 4.400 145.840 496.000 147.240 ;
        RECT 0.525 137.040 496.000 145.840 ;
        RECT 0.525 135.640 495.600 137.040 ;
        RECT 0.525 106.440 496.000 135.640 ;
        RECT 0.525 105.040 495.600 106.440 ;
        RECT 0.525 65.640 496.000 105.040 ;
        RECT 0.525 64.240 495.600 65.640 ;
        RECT 0.525 58.840 496.000 64.240 ;
        RECT 0.525 57.440 495.600 58.840 ;
        RECT 0.525 55.440 496.000 57.440 ;
        RECT 4.400 54.040 495.600 55.440 ;
        RECT 0.525 52.040 496.000 54.040 ;
        RECT 4.400 50.640 495.600 52.040 ;
        RECT 0.525 48.640 496.000 50.640 ;
        RECT 4.400 47.240 495.600 48.640 ;
        RECT 0.525 45.240 496.000 47.240 ;
        RECT 4.400 43.840 495.600 45.240 ;
        RECT 0.525 41.840 496.000 43.840 ;
        RECT 0.525 40.635 495.600 41.840 ;
  END
END fpga_top
END LIBRARY

